library verilog;
use verilog.vl_types.all;
entity DMem is
    port(
        DataOut         : out    vl_logic_vector(31 downto 0);
        DataAdr         : in     vl_logic_vector(7 downto 0);
        DataIn          : in     vl_logic_vector(31 downto 0);
        DMemW           : in     vl_logic;
        DMemR           : in     vl_logic;
        clk             : in     vl_logic
    );
end DMem;
