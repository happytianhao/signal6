library verilog;
use verilog.vl_types.all;
entity Mips is
end Mips;
